use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
library work;
use work.common.all;
entity imem is
port(
addr : in std_logic_vector(5 downto 0);
dout : out word);
end imem;
architecture behavioral of imem is
type rom_arr is array(0 to 46) of word;
constant mem:rom_arr:=
(
x"00000737" ,--8 0000 37070000 lui a4,%hi(lfsr.2565) 0000 0000 0000 0000 0000 0111 0011 0111
x"00075503" ,--9 0004 03550700 lhu a0,%lo(lfsr.2565)(a4) 0000 0000 0000 0111 0101 0101 0000 0011
x"00000013", -- 0008 13000000 nop
x"00755793" ,--10 000c 93577500 srli a5,a0,7 0000 0000 0111 0101 0101 0111 1001 0011
x"00000013", -- 0010 13000000 nop
x"00F547B3" ,--11 0014 B347F500 xor a5,a0,a5 0000 0000 1111 0101 0100 0111 1011 0011
x"00000013", -- 0018 13000000 nop
x"00979513" ,--12 001c 13959700 slli a0,a5,9
x"00000013", -- 0020 13000000 nop
x"00F54533" ,--13 0024 3345F500 xor a0,a0,a5
x"00000013", -- 0028 13000000 nop
x"01051513", --14 002c 13150501 slli a0,a0,16
x"00000013", -- 0030 13000000 nop
x"01055513" ,--15 0034 13550501 srli a0,a0,16
x"00000013", -- 0038 13000000 nop
x"00D55793" ,--16 003c 9357D500 srli a5,a0,13
x"00000013", -- 0040 13000000 nop
x"00F54533" ,--17 0044 3345F500 xor a0,a0,a5
x"00000013", -- 0048 13000000 nop
x"00A71023" ,--18 004c 2310A700 sh a0,%lo(lfsr.2565)(a4) 0000 0000 1010 0111 0001 0000 0010 0011
x"00008067", --19 0050 67800000 ret 0000 0000 0000 0000 1000 0000 0110 0111
--20 .size lfsr3, .-lfsr3
--21 .align 2
--22 .globl main
--23 .type main, @function
--24 main:
x"FF010113" ,--25 0054 130101FF addi sp,sp,-16 1111 1111 0000 0001 0000 0001 0001 0011 sp=-16
x"00000013", -- 0060 13000000 nop
x"00112623" ,--26 0064 23261100 sw ra,12(sp) 0000 0000 0001 0001 0010 01100010 0011 ra= -4
x"00812423" ,--27 006c 23248100 sw s0,8(sp)s0=-8
x"00912223" ,--28 0074 23229100 sw s1,4(sp)s1=-12
x"00000437" ,--29 007c 37040000 lui s0,%hi(outputs)0000 0000 0000 0000 0000 0100 0011 0111
x"00000013", -- 0080 13000000 nop
x"00040413" ,--30 0084 13040400 addi s0,s0,%lo(outputs)
x"00000013", -- 0088 13000000 nop
x"01E40493" ,--31 008c 9304E401 addi s1,s0,30
--32 .L3:
x"00000013", -- 0089 13000000 nop
x"00000097" ,--33 0094 97000000 call lfsr3 0000 0000 1001 0111
x"00000013", -- 0098 13000000 nop
x"000080E7" ,--33 009c E7800000 0000 0000 0000 0000 1000 0000 1110 0111
x"00000013", -- 00a0 13000000 nop
x"00A40023" ,--34 0094 2300A400 sb a0,0(s0)
x"00000013", -- 0098 13000000 nop
x"00140413" ,--35 009c 13041400 addi s0,s0,1
x"00000013", -- 00a0 13000000 nop
x"FC940EE3" ,--36 00a4 E31894FE bne s0,s1,.L3 11111100100101000000111011100011--11100
x"00000513", --37 0060 13050000 li a0,0
x"00C12083" ,--38 0064 8320C100 lw ra,12(sp)
x"00812403" ,--39 0068 03248100 lw s0,8(sp)
x"00412483" ,--40 006c 83244100 lw s1,4(sp)
x"01010113" ,--41 0070 13010101 addi sp,sp,16
x"00008067");--42 0074 67800000 jr ra -
- 13000000 nop
--43 .size main, .-main
--44 .comm outputs,30,4
--45 .section .sdata,"aw"
--46 .align 1
-- 47 .type lfsr.2565, @object
-- 48 .size lfsr.2565, 2
--49 lfsr.2565:
--50 0000 E1AC .half -21279
--51 .ident "GCC: (GNU) 8.2.0"
begin
    dout<=mem(conv_integer(addr));
    end behavioral;